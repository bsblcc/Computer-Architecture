module arm_alu_adder (
    input [31:0] operand_a,
    input [31:0] operand_b,
    input carry_in,
    output [31:0] out,

);
endmodule