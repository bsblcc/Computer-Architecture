////
//// Internal signal constants
////
